* Qucs 0.0.19  /home/fx/Arduino_stm32/batteryTester3/schematics/qucs19/simple.sch

.SUBCKT NMOSFETs_IRLZ44N  gnd  _net2 _net1 _net3
MM1 _net9 _net7 _net8 _net8 MMOD_M1 L=100u W=100u 
.MODEL MMOD_M1 NMOS(Is=1e-32 Vt0=2.08819 Lambda=0.0038193 Kp=67.9211 Cgso=1.59143e-05 Cgdo=3.04562e-08 Gamma=0 Phi=0.6) 
RRS _net8 _net3 0.014066
DD1 _net3 _net1 DMOD_D1 
.MODEL DMOD_D1 D(Is=4.4574e-09 Rs=0.007275 N=1.40246 Bv=55 Ibv=0.00025 Eg=1.14011 Xti=3.00078 Tt=0 Cj0=8.92434e-10 Vj=4.94724 M=0.75496 Fc=0.5) 
RRDS _net3 _net1 2.2e+06
RRD _net9 _net1 0.00179971
RRG _net2 _net7 2.4114
DD2 _net4 _net5 DMOD_D2 
.MODEL DMOD_D2 D(Is=1e-32 N=50 Cj0=1.15401e-09 Vj=0.859156 M=0.642548 Fc=1e-08) 
DD3 gnd _net5 DMOD_D3 
.MODEL DMOD_D3 D(Is=1e-10 N=0.4 Rs=3e-06 M=0.5 Cj0=1e-14 Vj=0.7) 
RRL _net5 _net10 1
FFI2 _net7 _net9 VFI2 -1
VFI2 _net4 _cnet0 DC 0
VdcVFI2 _cnet0 gnd DC 0
EEV16 _net10 gnd _net9 _net7 1
CCAP _net11 _net10 3.64838e-09
FFI1 _net7 _net9 VFI1 -1
VFI1 _net11 _cnet1 DC 0
VdcVFI1 _cnet1 _net6 DC 0
RRCAP _net6 _net10 1
DD4 gnd _net6 DMOD_D4 
.MODEL DMOD_D4 D(Is=1e-10 N=0.4 M=0.5 Cj0=1e-14 Vj=0.7) 
.ENDS


.SUBCKT Ideal_OpAmp gnd in_p in_m out AOLDC=106 GBP=1e6 RO=75 VLIMP=14 VLIMN=-14 
.PARAM OLG = {10**(AOLDC/20)}
.PARAM Fg = {GBP/OLG}
.PARAM pi = 3.14159
.PARAM C1 = {1e-3/sqrt(2*pi*fg)}
.PARAM R1 = {1e3/sqrt(2*pi*fg)}
ESRC1 _net0 0 in_p in_m OLG
R2 out  _net1 RO
R1 nC  _net0 R1
C1 nC  0 C1
B1 _net1  0  V = V(nC)*u(VLIMP-V(nC))*u(V(nC)-VLIMN)+VLIMP*u(V(nC)-VLIMP)+VLIMN*u(VLIMN-V(nC)) 
.ENDS
           

V2 _net0 0 DC 4
XIRLZ44N 0  gate _net1 SHUNT NMOSFETs_IRLZ44N
R1 _net1 _net0  2
R2 0 SHUNT  0.1
R5 0 _net2  820
XOP4 0  SHUNT _net2 _net3 Ideal_OpAmp GBP=1E6 AOLDC=106 RO=75 VLIMP=3.3 VLIMN=0
R6 _net3 _net2  22K
XOP3 0  _net4 _net3 gate Ideal_OpAmp GBP=1E6 AOLDC=106 RO=75 VLIMP=3.3 VLIMN=0
V5 _net4 0 DC 0.1
.control
echo "" > spice4qucs.cir.noise
echo "" > spice4qucs.cir.pz
tran 5e-05 0.01 0 
write simple_tran.txt v(SHUNT) v(gate) 
destroy all
reset

exit
.endc
.END
